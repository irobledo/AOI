LIBRARY ieee;
USE ieee.STD_LOGIC_1164.all;
ENTITY gateNOTE IS
  PORT (
   e0,e1   : IN STD_LOGIC; 
   s       : OUT STD_LOGIC
       );
END gateNOTE;
