ARCHITECTURE flujo OF gateNOTE IS
-- Parte declarativa

BEGIN
-- Descripci�n de la arquitectura

 s<= e0 OR e1;

END flujo;

----------------------------------------------------------------------

