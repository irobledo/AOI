LIBRARY ieee;
USE ieee.STD_LOGIC_1164.all;
ENTITY gateOR2 IS
  PORT (
   e0,e1   : IN STD_LOGIC; 
   s       : OUT STD_LOGIC
       );
END gateOR2;
